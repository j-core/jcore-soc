library ieee;
use ieee.std_logic_1164.all;
use std.textio.all;
use ieee.std_logic_textio.all;
use ieee.numeric_std.all;

use work.cache_pack.all;
use work.cpu2j0_pack.all;
use work.data_bus_pack.all;
use work.dma_pack.all;

entity dcache_tb is
end dcache_tb;

-- dhrystone special tb
--   acc_vect 72 bits (normal vector 68 bits) entexsion is en bit
--   acc_vect includes cpu en=0 cycle
--   dhrystone loop control in vector

architecture tb of dcache_tb is

type acc_vect_t is array (0 to 2047)  of std_logic_vector( 71 downto 0);
type ddr_ram_t  is array (0 to 2**14-1)  of std_logic_vector( 31 downto 0);

   signal rst   : std_logic;
   signal rst_46nsdel   : std_logic;
   signal clk125   : std_logic;
   signal clk200   : std_logic;

   signal a0     : cpu_data_o_t;
   signal y0     : cpu_data_i_t;
   signal sa0    : dcache_snoop_io_t;
   signal sy0    : dcache_snoop_io_t;
   signal sy0_1del : dcache_snoop_io_t;
   signal ra0    : dcache_ram_o_t;
   signal ry0    : dcache_ram_i_t;
   signal ma0    : mem_i_t;
   signal my0    : mem_o_t;

   signal a1     : cpu_data_o_t;
   signal y1     : cpu_data_i_t;
   signal ra1    : dcache_ram_o_t;
   signal ry1    : dcache_ram_i_t;
   signal ma1    : mem_i_t;
   signal my1    : mem_o_t;

   signal ma    : mem_i_t;
   signal my    : mem_o_t;

   signal  m1_o   : cpu_data_i_t;
   signal  m1_i   : cpu_data_o_t;
   signal  m2_o   : bus_ddr_i_t;
   signal  m2_i   : bus_ddr_o_t;
   signal  mem_o : cpu_data_o_t;
   signal  mem_i : cpu_data_i_t;

   signal ctrl  : cache_ctrl_t;
   signal my_1delay : mem_o_t;
   signal ma_rdy_1wait_sig : std_logic;

   signal cavec  : std_logic_vector( 67 downto 0 );

   signal acc_vect : acc_vect_t;
   signal ddr_ram  : ddr_ram_t := ( others => x"A5A5A5A5" );
   signal acksp_pointer_thisc : std_logic_vector(10 downto 0);
   signal acksp_pointer_thisr : std_logic_vector(10 downto 0);
   signal mis_counter_thisc : std_logic_vector(10 downto 0);
   signal mis_counter_thisr : std_logic_vector(10 downto 0);
   signal y_ack_1del_thisc : std_logic;
   signal y_ack_1del_thisr : std_logic;
   signal observe_dcache_waitsig  : std_logic;

   for mem0 : dcache_ram
     use configuration work.dcache_ram_infer;
   for mem1 : dcache_ram
     use configuration work.dcache_ram_infer;

begin

  --
  rst <= '1', '0' after 15 ns;
  rst_46nsdel <= rst after 46 ns;
  clk125 <= '0' after 4   ns when clk125 = '1' else '1' after 4   ns;
  clk200 <= '0' after 2.5 ns when clk200 = '1' else '1' after 2.5 ns;

-- .+....1....+....1....+....1....+....1....+....1....+....1....+....1....+....1
  dut0 : dcache     port map ( rst => rst,
    clk125 => clk125, clk200 => clk200, a => a0,
    lock => '0',      y => y0,          sa => sa0,
    sy => sy0,        ra => ra0,        ry => ry0,
    ma => ma0,        my => my0 ,       ctrl   => ctrl );
  mem0 : dcache_ram      port map ( rst => rst,
    clk125 => clk125,
    clk200 => clk200, ra => ry0, ry => ra0 );

  dut1 : dcache     port map ( rst => rst,
    clk125 => clk125, clk200 => clk200, a => a1,
    lock => '0',      y => y1,          sa => sy0,
    sy => sa0,        ra => ra1,        ry => ry1,
    ma => ma1,        my => my1 ,       ctrl   => ctrl );
  mem1 : dcache_ram      port map ( rst => rst,
    clk125 => clk125,
    clk200 => clk200, ra => ry1, ry => ra1 );

  dut2 : bus_mux_typeb port map (
    clk    => clk200, 
    rst    => rst, 
    m1_o   => m1_o,
    m1_i   => m1_i,
    m2_o   => m2_o,
    m2_i   => m2_i,
    mem_o  => mem_o,
    mem_i  => mem_i);

  -- connection around bus_mux_typeb
  m1_i.en <= my0.en;
  m1_i.a  <= x"0" & my0.a;
  m1_i.wr <= my0.wr;
  m1_i.we <= my0.we;
  m1_i.d  <= my0.d ;
  m1_i.rd <= my0.en and (not my0.wr);
  ma0.ack <= m1_o.ack;
  ma0.d   <= m1_o.d  ;

  m2_i.en <= my1.en;
  m2_i.a  <= x"0" & my1.a;
  m2_i.wr <= my1.wr;
  m2_i.we <= my1.we;
  m2_i.d  <= my1.d ;
  ma1.ack <= m2_o.ack;
  ma1.d   <= m2_o.d  ;

  my.en   <= mem_o.en;
  my.a    <= mem_o.a(27 downto 0);
  my.wr   <= mem_o.wr;
  my.we   <= mem_o.we;
  my.d    <= mem_o.d ;
  mem_i.ack <= ma.ack;
  mem_i.d   <= ma.d;

  sy0_1del <= sy0 after 8 ns;

-- .+....1....+....1....+....1....+....1....+....1....+....1....+....1....+....1
--  sa.en <= '0';
--  sa.al <= (others => '0');
-- .+....1....+....1....+....1....+....1....+....1....+....1....+....1....+....1
  -- cache on/off selection
  -- --------------------------------------------------------------------------
    ctrl.en  <= '1' ; -- cache on
--  ctrl.en  <= '0' ; -- cache off
-- --------------------------------------------------------------------------
    ctrl.inv <= '0' ; -- no invalidate 
-- --------------------------------------------------------------------------

--  valid_rest : process( acksp_pointer_thisr, y_ack_1del_thisr, rst_46nsdel)
--  begin
--    if(y_ack_1del_thisr = '1') and
--      (acksp_pointer_thisr(2 downto 0) = b"111") then
--      a.a  <= x"0aaaaaa0";
--      a.en <= '0';
--      a.wr <= '0';
--      a.we <= x"0";
--      a.d  <= x"00000000";
--    else
      a0.a  <= x"0" &
               acc_vect(vtoi(acksp_pointer_thisr))(59 downto 32);
      a0.en <= acc_vect(vtoi(acksp_pointer_thisr))(68) and
               (not acc_vect(vtoi(acksp_pointer_thisr))(69));
      a0.wr <= acc_vect(vtoi(acksp_pointer_thisr))(64) and
               (not acc_vect(vtoi(acksp_pointer_thisr))(69));
      a0.we <= acc_vect(vtoi(acksp_pointer_thisr))(63 downto 60);
      a0.d  <= acc_vect(vtoi(acksp_pointer_thisr))(31 downto  0);

      a1.a  <= x"0" &
               acc_vect(vtoi(acksp_pointer_thisr))(59 downto 32);
      a1.en <= acc_vect(vtoi(acksp_pointer_thisr))(68) and
               acc_vect(vtoi(acksp_pointer_thisr))(69);
      a1.wr <= acc_vect(vtoi(acksp_pointer_thisr))(64) and
               acc_vect(vtoi(acksp_pointer_thisr))(69);
      a1.we <= acc_vect(vtoi(acksp_pointer_thisr))(63 downto 60);
      a1.d  <= acc_vect(vtoi(acksp_pointer_thisr))(31 downto  0);
--    end if;
--  end process;

  ma.d <= (ddr_ram(vtoi(my.a(15 downto 2)))) and
   (
    ma.ack & ma.ack & ma.ack & ma.ack &
    ma.ack & ma.ack & ma.ack & ma.ack &
    ma.ack & ma.ack & ma.ack & ma.ack &
    ma.ack & ma.ack & ma.ack & ma.ack &
    ma.ack & ma.ack & ma.ack & ma.ack &
    ma.ack & ma.ack & ma.ack & ma.ack &
    ma.ack & ma.ack & ma.ack & ma.ack &
    ma.ack & ma.ack & ma.ack & ma.ack 
   ) ;

  my_1delay <= my after 5 ns;

  -- --------------------------------------------------------------------------
  gen_ready_1wait : process (my, my_1delay)
    variable mem_rdy_1wait : std_logic;
  begin
    if (my_1delay.en = '1') and
       (my.en        = '1') and
       (my_1delay.a = my.a) then mem_rdy_1wait := '1';
     else                        mem_rdy_1wait := '0';
     end if;
     ma_rdy_1wait_sig <=     mem_rdy_1wait;
  end process;
  -- --------------------------------------------------------------------------
  -- 1 wait
  ma.ack <= ma_rdy_1wait_sig;
  -- --------------------------------------------------------------------------
  -- 0 wait
--  ma.ack <= my.en;
  -- --------------------------------------------------------------------------
  observe_dcache_waitsig <= a0.en and (not y0.ack);

  ackfsm : process(acksp_pointer_thisr, mis_counter_thisr, y_ack_1del_thisr,
     y0.ack, y1.ack, my.av, ma.ack , a0.en, a1.en, rst, rst_46nsdel )
   variable acksp_pointer_this : std_logic_vector(10 downto 0);
   variable mis_counter_this : std_logic_vector(10 downto 0);
   variable y_ack_1del_this  : std_logic;
  begin
   acksp_pointer_this := acksp_pointer_thisr;
   mis_counter_this := mis_counter_thisr;
   y_ack_1del_this  := y_ack_1del_thisr;

   if(rst = '1') or (rst_46nsdel /= '0') then
        -- acksp_pointer_this update disabled
   elsif(y0.ack = '1') or (y1.ack = '1') or
        ((a0.en = '0') and (a1.en = '0')) then
     acksp_pointer_this := std_logic_vector(unsigned(acksp_pointer_this) + 1);
     -- dhrystone loop control
     if (acksp_pointer_this = b"101" & x"5b") then -- 0x55b (dec 1371)
       acksp_pointer_this :=  b"001" & x"8a";      -- 0x18a (dec  394)
     end if;
   end if;
   if((my.av = '1') and (ma.ack = '1')) then
     mis_counter_this := std_logic_vector(unsigned(mis_counter_this) + 1);
   end if;
   y_ack_1del_this := (y0.ack or y1.ack);

   acksp_pointer_thisc <= acksp_pointer_this;
   mis_counter_thisc <= mis_counter_this;
   y_ack_1del_thisc  <= y_ack_1del_this ;
  end process;

  p0_r0_125fsm : process(clk125, rst)
  begin
     if rst = '1' then
        acksp_pointer_thisr <= b"000" & x"00";
        y_ack_1del_thisr  <= '0';
     elsif clk125 = '1' and clk125'event then
        acksp_pointer_thisr <= acksp_pointer_thisc;
        y_ack_1del_thisr  <= y_ack_1del_thisc ;
     end if;
  end process;

  p0_r0_200fsm : process(clk200, rst)
  begin
     if rst = '1' then
        mis_counter_thisr <= b"000" & x"00";
     elsif clk200 = '1' and clk200'event then
        mis_counter_thisr <= mis_counter_thisc;
     end if;
  end process;

  ddr_raminit : process(rst, my)
  begin
   if rst = '1' then
   ddr_ram(    0) <= x"000000cc";
   ddr_ram(    1) <= x"00000000";
   ddr_ram(   61) <= x"000097fc";
   ddr_ram(   62) <= x"00009ffc";
   ddr_ram(   63) <= x"00000288";
   ddr_ram(   76) <= x"0000c450";
   ddr_ram(   77) <= x"0000c44c";
   ddr_ram(   89) <= x"0000c454";
   ddr_ram(   90) <= x"0000c44c";
   ddr_ram(   91) <= x"00000894";
   ddr_ram(  139) <= x"0000c454";
   ddr_ram(  140) <= x"00000138";
   ddr_ram(  141) <= x"000009c0";
   ddr_ram(  142) <= x"00000894";
   ddr_ram(  151) <= x"0000c520";
   ddr_ram(  152) <= x"0000c450";
   ddr_ram(  153) <= x"0000c451";
   ddr_ram(  160) <= x"0000c450";
   ddr_ram(  161) <= x"0000c520";
   ddr_ram(  198) <= x"00000384";
   ddr_ram(  288) <= x"4e470009";
   ddr_ram(  289) <= x"000031e8";
   ddr_ram(  290) <= x"0000c448";
   ddr_ram(  291) <= x"0000c454";
   ddr_ram(  292) <= x"44485259";
   ddr_ram(  293) <= x"53544f4e";
   ddr_ram(  294) <= x"45205052";
   ddr_ram(  295) <= x"4f475241";
   ddr_ram(  296) <= x"4d2c2053";
   ddr_ram(  297) <= x"4f4d4520";
   ddr_ram(  298) <= x"53545249";
   ddr_ram(  299) <= x"4d2c2031";
   ddr_ram(  300) <= x"27535420";
   ddr_ram(  301) <= x"0000a370";
   ddr_ram(  316) <= x"00000268";
   ddr_ram(  317) <= x"0000023c";
   ddr_ram(  318) <= x"4d2c2032";
   ddr_ram(  319) <= x"274e4420";
   ddr_ram(  320) <= x"00000944";
   ddr_ram(  321) <= x"0000c520";
   ddr_ram(  322) <= x"00000894";
   ddr_ram(  323) <= x"0000c458";
   ddr_ram(  324) <= x"00009d34";
   ddr_ram(  325) <= x"000008a4";
   ddr_ram(  326) <= x"00000170";
   ddr_ram(  327) <= x"0000c451";
   ddr_ram(  328) <= x"4d2c2033";
   ddr_ram(  329) <= x"00000924";
   ddr_ram(  486) <= x"00001acc";
   ddr_ram(  487) <= x"00000110";
   ddr_ram(  583) <= x"00c80fa0";
   ddr_ram(  584) <= x"0000c44c";
   ddr_ram(  617) <= x"00000924";
   ddr_ram(  618) <= x"00002d14";
   ddr_ram(  636) <= x"000009b0";
   ddr_ram(  637) <= x"00002630";
   ddr_ram( 3184) <= x"000035e4";
   ddr_ram( 3185) <= x"0000322c";
   ddr_ram( 3186) <= x"000035e4";
   ddr_ram( 3207) <= x"000030e4";
   ddr_ram( 3208) <= x"00007ae8";
   ddr_ram( 3209) <= x"00009cb8";
   ddr_ram( 7866) <= x"00007be8";
   ddr_ram( 7894) <= x"4e470000";
   ddr_ram( 7930) <= x"00000100";
   ddr_ram(10210) <= x"00000000";
   ddr_ram(10219) <= x"4e474e47";
   ddr_ram(10227) <= x"4e474e47";
   ddr_ram(12564) <= x"41420000";
   elsif (my.en = '1') and (my.wr = '1') then
     for i in 0 to 3 loop
       if(my.we(i) = '1') then
         ddr_ram(vtoi(my.a(15 downto 2)))(8 * i + 7 downto 8 * i)
         <= my.d                         (8 * i + 7 downto 8 * i);
       end if;
     end loop;
   end if;
   end process;

-- ---- cpu access dump ------
  process
    file f0 : text is out "cpu0.acc";
    variable l : line;
  begin

    wait for 1 ns;
    if(y0.ack = '1') then
      hwrite(     l, a0.a );   write(l, string'(" "));
      if(a0.wr = '1') then
           hwrite(l, a0.d );   write(l, string'(" "));
      else hwrite(l, y0.d );   write(l, string'(" "));
      end if;
       write(     l, a0.wr );  write(l, string'(" "));
      -- write line --------------
      writeline(f0, l);
      deallocate(l);
    end if;
    wait for 7 ns;
  end process;

-- ---- bus write dump ------
  process
    file f1 : text is out "bus.acc";
    variable l1 : line;
  begin

    wait for 1 ns;
    if(ma.ack = '1') and (my.wr = '1') then
      hwrite(l1, my.a );   write(l1, string'(" "));
      hwrite(l1, my.d );   write(l1, string'(" "));
      -- write line --------------
      writeline(f1, l1);
      deallocate(l1);
    end if;
    wait for 4 ns;
  end process;

-- ---- snoop write dump (en and next cycle) ------
  process
    file f2 : text is out "snoopo.acc";
    variable l2 : line;
  begin

    wait for 1 ns;
    if(sy0.en = '1') or (sy0_1del.en = '1') then
      hwrite(l2, sy0.al & '0' );
      -- write line --------------
      writeline(f2, l2);
      deallocate(l2);
    end if;
    wait for 7 ns;
  end process;

-- ---- snoop write dump ------
    



  -- vector           eww
  --                  nre  adr    data
  --                  ||||_____||______|
  -- prepare hit entry
  --
-- cpu_sim load/store vector
-- initialize finish
  acc_vect(   0) <= x"000000000000000000";
  acc_vect(   1) <= x"000000000000000000";
  acc_vect(   2) <= x"000000000000000000";
  acc_vect(   3) <= x"1000000000000000CC";
  acc_vect(   4) <= x"100000000400000000";
  acc_vect(   5) <= x"000000000000000000";
  acc_vect(   6) <= x"000000000000000000";
  acc_vect(   7) <= x"000000000000000000";
  acc_vect(   8) <= x"000000000000000000";
  acc_vect(   9) <= x"000000000000000000";
  acc_vect(  10) <= x"000000000000000000";
  acc_vect(  11) <= x"000000000000000000";
  acc_vect(  12) <= x"000000000000000000";
  acc_vect(  13) <= x"000000000000000000";
  acc_vect(  14) <= x"000000000000000000";
  acc_vect(  15) <= x"000000000000000000";
  acc_vect(  16) <= x"000000000000000000";
  acc_vect(  17) <= x"000000000000000000";
  acc_vect(  18) <= x"000000000000000000";
  acc_vect(  19) <= x"000000000000000000";
  acc_vect(  20) <= x"000000000000000000";
  acc_vect(  21) <= x"000000000000000000";
  acc_vect(  22) <= x"10000000F4000097FC";
  acc_vect(  23) <= x"10000000F800009FFC";
  acc_vect(  24) <= x"10000000FC00000288";
  acc_vect(  25) <= x"000000000000000000";
  acc_vect(  26) <= x"000000000000000000";
  acc_vect(  27) <= x"000000000000000000";
  acc_vect(  28) <= x"000000000000000000";
  acc_vect(  29) <= x"11F0009FF800000000";
  acc_vect(  30) <= x"11F0009FF400000000";
  acc_vect(  31) <= x"11F0009FF000000000";
  acc_vect(  32) <= x"11F0009FEC00000000";
  acc_vect(  33) <= x"11F0009FE800000000";
  acc_vect(  34) <= x"11F0009FE400000000";
  acc_vect(  35) <= x"11F0009FE0000097FC";
  acc_vect(  36) <= x"11F0009FDC000000F2";
  acc_vect(  37) <= x"000000000000000000";
  acc_vect(  38) <= x"000000000000000000";
  acc_vect(  39) <= x"1000000484000031E8";
  acc_vect(  40) <= x"000000000000000000";
  acc_vect(  41) <= x"000000000000000000";
  acc_vect(  42) <= x"000000000000000000";
  acc_vect(  43) <= x"000000000000000000";
  acc_vect(  44) <= x"11F0009F8000009F84";
  acc_vect(  45) <= x"000000000000000000";
  acc_vect(  46) <= x"11F0009F7C000002A2";
  acc_vect(  47) <= x"000000000000000000";
  acc_vect(  48) <= x"000000000000000000";
  acc_vect(  49) <= x"000000000000000000";
  acc_vect(  50) <= x"000000000000000000";
  acc_vect(  51) <= x"000000000000000000";
  acc_vect(  52) <= x"100000321C000030E4";
  acc_vect(  53) <= x"100000322000007AE8";
  acc_vect(  54) <= x"100000322400009CB8";
  acc_vect(  55) <= x"000000000000000000";
  acc_vect(  56) <= x"000000000000000000";
  acc_vect(  57) <= x"000000000000000000";
  acc_vect(  58) <= x"11F0009F7800000000";
  acc_vect(  59) <= x"000000000000000000";
  acc_vect(  60) <= x"11F0009F74000031E8";
  acc_vect(  61) <= x"000000000000000000";
  acc_vect(  62) <= x"11F0009F7000000000";
  acc_vect(  63) <= x"000000000000000000";
  acc_vect(  64) <= x"11F0009F6C00000000";
  acc_vect(  65) <= x"11F0009F6800000000";
  acc_vect(  66) <= x"11F0009F6400009F7C";
  acc_vect(  67) <= x"11F0009F6000003202";
  acc_vect(  68) <= x"10000031C0000035E4";
  acc_vect(  69) <= x"000000000000000000";
  acc_vect(  70) <= x"000000000000000000";
  acc_vect(  71) <= x"11F0009F5C00000034";
  acc_vect(  72) <= x"000000000000000000";
  acc_vect(  73) <= x"000000000000000000";
  acc_vect(  74) <= x"000000000000000000";
  acc_vect(  75) <= x"11F0009F5800009F5C";
  acc_vect(  76) <= x"000000000000000000";
  acc_vect(  77) <= x"000000000000000000";
  acc_vect(  78) <= x"000000000000000000";
  acc_vect(  79) <= x"000000000000000000";
  acc_vect(  80) <= x"000000000000000000";
  acc_vect(  81) <= x"000000000000000000";
  acc_vect(  82) <= x"1000009F5800009F5C";
  acc_vect(  83) <= x"10000031C40000322C";
  acc_vect(  84) <= x"000000000000000000";
  acc_vect(  85) <= x"000000000000000000";
  acc_vect(  86) <= x"000000000000000000";
  acc_vect(  87) <= x"000000000000000000";
  acc_vect(  88) <= x"1000009F5C00000034";
  acc_vect(  89) <= x"000000000000000000";
  acc_vect(  90) <= x"11F0009F5800009F5C";
  acc_vect(  91) <= x"000000000000000000";
  acc_vect(  92) <= x"000000000000000000";
  acc_vect(  93) <= x"000000000000000000";
  acc_vect(  94) <= x"000000000000000000";
  acc_vect(  95) <= x"000000000000000000";
  acc_vect(  96) <= x"000000000000000000";
  acc_vect(  97) <= x"000000000000000000";
  acc_vect(  98) <= x"000000000000000000";
  acc_vect(  99) <= x"000000000000000000";
  acc_vect( 100) <= x"1000007AE800007BE8";
  acc_vect( 101) <= x"000000000000000000";
  acc_vect( 102) <= x"000000000000000000";
  acc_vect( 103) <= x"000000000000000000";
  acc_vect( 104) <= x"000000000000000000";
  acc_vect( 105) <= x"000000000000000000";
  acc_vect( 106) <= x"1000007BE800000100";
  acc_vect( 107) <= x"000000000000000000";
  acc_vect( 108) <= x"000000000000000000";
  acc_vect( 109) <= x"000000000000000000";
  acc_vect( 110) <= x"000000000000000000";
  acc_vect( 111) <= x"000000000000000000";
  acc_vect( 112) <= x"000000000000000000";
  acc_vect( 113) <= x"000000000000000000";
  acc_vect( 114) <= x"000000000000000000";
  acc_vect( 115) <= x"000000000000000000";
  acc_vect( 116) <= x"000000000000000000";
  acc_vect( 117) <= x"000000000000000000";
  acc_vect( 118) <= x"000000000000000000";
  acc_vect( 119) <= x"11F0007BE8000000CC";
  acc_vect( 120) <= x"000000000000000000";
  acc_vect( 121) <= x"000000000000000000";
  acc_vect( 122) <= x"000000000000000000";
  acc_vect( 123) <= x"11F0009F5C00000034";
  acc_vect( 124) <= x"000000000000000000";
  acc_vect( 125) <= x"000000000000000000";
  acc_vect( 126) <= x"000000000000000000";
  acc_vect( 127) <= x"000000000000000000";
  acc_vect( 128) <= x"1000009F5800009F5C";
  acc_vect( 129) <= x"000000000000000000";
  acc_vect( 130) <= x"10000031C8000035E4";
  acc_vect( 131) <= x"000000000000000000";
  acc_vect( 132) <= x"000000000000000000";
  acc_vect( 133) <= x"000000000000000000";
  acc_vect( 134) <= x"000000000000000000";
  acc_vect( 135) <= x"11F0009F5800009F5C";
  acc_vect( 136) <= x"000000000000000000";
  acc_vect( 137) <= x"000000000000000000";
  acc_vect( 138) <= x"000000000000000000";
  acc_vect( 139) <= x"000000000000000000";
  acc_vect( 140) <= x"000000000000000000";
  acc_vect( 141) <= x"000000000000000000";
  acc_vect( 142) <= x"1000009F5800009F5C";
  acc_vect( 143) <= x"000000000000000000";
  acc_vect( 144) <= x"000000000000000000";
  acc_vect( 145) <= x"000000000000000000";
  acc_vect( 146) <= x"1000009F5C00000034";
  acc_vect( 147) <= x"000000000000000000";
  acc_vect( 148) <= x"000000000000000000";
  acc_vect( 149) <= x"000000000000000000";
  acc_vect( 150) <= x"000000000000000000";
  acc_vect( 151) <= x"11F0007AF400000034";
  acc_vect( 152) <= x"000000000000000000";
  acc_vect( 153) <= x"000000000000000000";
  acc_vect( 154) <= x"1000009F6000003202";
  acc_vect( 155) <= x"000000000000000000";
  acc_vect( 156) <= x"000000000000000000";
  acc_vect( 157) <= x"1000009F6400009F7C";
  acc_vect( 158) <= x"000000000000000000";
  acc_vect( 159) <= x"1000009F6800000000";
  acc_vect( 160) <= x"000000000000000000";
  acc_vect( 161) <= x"1000009F6C00000000";
  acc_vect( 162) <= x"000000000000000000";
  acc_vect( 163) <= x"1000009F7000000000";
  acc_vect( 164) <= x"000000000000000000";
  acc_vect( 165) <= x"1000009F74000031E8";
  acc_vect( 166) <= x"000000000000000000";
  acc_vect( 167) <= x"000000000000000000";
  acc_vect( 168) <= x"000000000000000000";
  acc_vect( 169) <= x"1000009F7800000000";
  acc_vect( 170) <= x"000000000000000000";
  acc_vect( 171) <= x"000000000000000000";
  acc_vect( 172) <= x"000000000000000000";
  acc_vect( 173) <= x"000000000000000000";
  acc_vect( 174) <= x"000000000000000000";
  acc_vect( 175) <= x"1000009F7C000002A2";
  acc_vect( 176) <= x"000000000000000000";
  acc_vect( 177) <= x"000000000000000000";
  acc_vect( 178) <= x"000000000000000000";
  acc_vect( 179) <= x"000000000000000000";
  acc_vect( 180) <= x"1000009F8000009F84";
  acc_vect( 181) <= x"10000004880000C448";
  acc_vect( 182) <= x"000000000000000000";
  acc_vect( 183) <= x"11F000C44800007AF8";
  acc_vect( 184) <= x"000000000000000000";
  acc_vect( 185) <= x"000000000000000000";
  acc_vect( 186) <= x"000000000000000000";
  acc_vect( 187) <= x"11F0009F8000009F84";
  acc_vect( 188) <= x"000000000000000000";
  acc_vect( 189) <= x"11F0009F7C000002AA";
  acc_vect( 190) <= x"000000000000000000";
  acc_vect( 191) <= x"000000000000000000";
  acc_vect( 192) <= x"000000000000000000";
  acc_vect( 193) <= x"000000000000000000";
  acc_vect( 194) <= x"000000000000000000";
  acc_vect( 195) <= x"100000321C000030E4";
  acc_vect( 196) <= x"100000322000007AE8";
  acc_vect( 197) <= x"100000322400009CB8";
  acc_vect( 198) <= x"000000000000000000";
  acc_vect( 199) <= x"000000000000000000";
  acc_vect( 200) <= x"000000000000000000";
  acc_vect( 201) <= x"11F0009F780000C448";
  acc_vect( 202) <= x"000000000000000000";
  acc_vect( 203) <= x"11F0009F74000031E8";
  acc_vect( 204) <= x"000000000000000000";
  acc_vect( 205) <= x"11F0009F7000000000";
  acc_vect( 206) <= x"000000000000000000";
  acc_vect( 207) <= x"11F0009F6C00000000";
  acc_vect( 208) <= x"11F0009F6800000000";
  acc_vect( 209) <= x"11F0009F6400009F7C";
  acc_vect( 210) <= x"11F0009F6000003202";
  acc_vect( 211) <= x"10000031C0000035E4";
  acc_vect( 212) <= x"000000000000000000";
  acc_vect( 213) <= x"000000000000000000";
  acc_vect( 214) <= x"11F0009F5C00000034";
  acc_vect( 215) <= x"000000000000000000";
  acc_vect( 216) <= x"000000000000000000";
  acc_vect( 217) <= x"000000000000000000";
  acc_vect( 218) <= x"11F0009F5800009F5C";
  acc_vect( 219) <= x"000000000000000000";
  acc_vect( 220) <= x"000000000000000000";
  acc_vect( 221) <= x"000000000000000000";
  acc_vect( 222) <= x"000000000000000000";
  acc_vect( 223) <= x"000000000000000000";
  acc_vect( 224) <= x"000000000000000000";
  acc_vect( 225) <= x"1000009F5800009F5C";
  acc_vect( 226) <= x"10000031C40000322C";
  acc_vect( 227) <= x"000000000000000000";
  acc_vect( 228) <= x"000000000000000000";
  acc_vect( 229) <= x"000000000000000000";
  acc_vect( 230) <= x"000000000000000000";
  acc_vect( 231) <= x"1000009F5C00000034";
  acc_vect( 232) <= x"000000000000000000";
  acc_vect( 233) <= x"11F0009F5800009F5C";
  acc_vect( 234) <= x"000000000000000000";
  acc_vect( 235) <= x"000000000000000000";
  acc_vect( 236) <= x"000000000000000000";
  acc_vect( 237) <= x"000000000000000000";
  acc_vect( 238) <= x"000000000000000000";
  acc_vect( 239) <= x"000000000000000000";
  acc_vect( 240) <= x"000000000000000000";
  acc_vect( 241) <= x"000000000000000000";
  acc_vect( 242) <= x"000000000000000000";
  acc_vect( 243) <= x"1000007AE800007BE8";
  acc_vect( 244) <= x"000000000000000000";
  acc_vect( 245) <= x"000000000000000000";
  acc_vect( 246) <= x"000000000000000000";
  acc_vect( 247) <= x"000000000000000000";
  acc_vect( 248) <= x"000000000000000000";
  acc_vect( 249) <= x"1000007BE8000000CC";
  acc_vect( 250) <= x"000000000000000000";
  acc_vect( 251) <= x"000000000000000000";
  acc_vect( 252) <= x"000000000000000000";
  acc_vect( 253) <= x"000000000000000000";
  acc_vect( 254) <= x"000000000000000000";
  acc_vect( 255) <= x"000000000000000000";
  acc_vect( 256) <= x"000000000000000000";
  acc_vect( 257) <= x"000000000000000000";
  acc_vect( 258) <= x"000000000000000000";
  acc_vect( 259) <= x"000000000000000000";
  acc_vect( 260) <= x"000000000000000000";
  acc_vect( 261) <= x"000000000000000000";
  acc_vect( 262) <= x"11F0007BE800000098";
  acc_vect( 263) <= x"000000000000000000";
  acc_vect( 264) <= x"000000000000000000";
  acc_vect( 265) <= x"000000000000000000";
  acc_vect( 266) <= x"11F0009F5C00000034";
  acc_vect( 267) <= x"000000000000000000";
  acc_vect( 268) <= x"000000000000000000";
  acc_vect( 269) <= x"000000000000000000";
  acc_vect( 270) <= x"000000000000000000";
  acc_vect( 271) <= x"1000009F5800009F5C";
  acc_vect( 272) <= x"000000000000000000";
  acc_vect( 273) <= x"10000031C8000035E4";
  acc_vect( 274) <= x"000000000000000000";
  acc_vect( 275) <= x"000000000000000000";
  acc_vect( 276) <= x"000000000000000000";
  acc_vect( 277) <= x"000000000000000000";
  acc_vect( 278) <= x"11F0009F5800009F5C";
  acc_vect( 279) <= x"000000000000000000";
  acc_vect( 280) <= x"000000000000000000";
  acc_vect( 281) <= x"000000000000000000";
  acc_vect( 282) <= x"000000000000000000";
  acc_vect( 283) <= x"000000000000000000";
  acc_vect( 284) <= x"000000000000000000";
  acc_vect( 285) <= x"1000009F5800009F5C";
  acc_vect( 286) <= x"000000000000000000";
  acc_vect( 287) <= x"000000000000000000";
  acc_vect( 288) <= x"000000000000000000";
  acc_vect( 289) <= x"1000009F5C00000034";
  acc_vect( 290) <= x"000000000000000000";
  acc_vect( 291) <= x"000000000000000000";
  acc_vect( 292) <= x"000000000000000000";
  acc_vect( 293) <= x"000000000000000000";
  acc_vect( 294) <= x"11F0007B2800000034";
  acc_vect( 295) <= x"000000000000000000";
  acc_vect( 296) <= x"000000000000000000";
  acc_vect( 297) <= x"1000009F6000003202";
  acc_vect( 298) <= x"000000000000000000";
  acc_vect( 299) <= x"000000000000000000";
  acc_vect( 300) <= x"1000009F6400009F7C";
  acc_vect( 301) <= x"000000000000000000";
  acc_vect( 302) <= x"1000009F6800000000";
  acc_vect( 303) <= x"000000000000000000";
  acc_vect( 304) <= x"1000009F6C00000000";
  acc_vect( 305) <= x"000000000000000000";
  acc_vect( 306) <= x"1000009F7000000000";
  acc_vect( 307) <= x"000000000000000000";
  acc_vect( 308) <= x"1000009F74000031E8";
  acc_vect( 309) <= x"000000000000000000";
  acc_vect( 310) <= x"000000000000000000";
  acc_vect( 311) <= x"000000000000000000";
  acc_vect( 312) <= x"1000009F780000C448";
  acc_vect( 313) <= x"000000000000000000";
  acc_vect( 314) <= x"000000000000000000";
  acc_vect( 315) <= x"000000000000000000";
  acc_vect( 316) <= x"000000000000000000";
  acc_vect( 317) <= x"000000000000000000";
  acc_vect( 318) <= x"1000009F7C000002AA";
  acc_vect( 319) <= x"000000000000000000";
  acc_vect( 320) <= x"000000000000000000";
  acc_vect( 321) <= x"000000000000000000";
  acc_vect( 322) <= x"000000000000000000";
  acc_vect( 323) <= x"1000009F8000009F84";
  acc_vect( 324) <= x"100000048C0000C454";
  acc_vect( 325) <= x"000000000000000000";
  acc_vect( 326) <= x"11F000C45400007B2C";
  acc_vect( 327) <= x"100000C44800007AF8";
  acc_vect( 328) <= x"000000000000000000";
  acc_vect( 329) <= x"11F0007B2C00007AF8";
  acc_vect( 330) <= x"100000C45400007B2C";
  acc_vect( 331) <= x"000000000000000000";
  acc_vect( 332) <= x"11F0007B3000000000";
  acc_vect( 333) <= x"000000000000000000";
  acc_vect( 334) <= x"11F0007B3400000002";
  acc_vect( 335) <= x"000000000000000000";
  acc_vect( 336) <= x"11F0007B3800000028";
  acc_vect( 337) <= x"100000049044485259";
  acc_vect( 338) <= x"000000000000000000";
  acc_vect( 339) <= x"11F0007B3C44485259";
  acc_vect( 340) <= x"100000049453544F4E";
  acc_vect( 341) <= x"000000000000000000";
  acc_vect( 342) <= x"11F0007B4053544F4E";
  acc_vect( 343) <= x"100000049845205052";
  acc_vect( 344) <= x"000000000000000000";
  acc_vect( 345) <= x"11F0007B4445205052";
  acc_vect( 346) <= x"100000049C4F475241";
  acc_vect( 347) <= x"000000000000000000";
  acc_vect( 348) <= x"11F0007B484F475241";
  acc_vect( 349) <= x"10000004A04D2C2053";
  acc_vect( 350) <= x"000000000000000000";
  acc_vect( 351) <= x"11F0007B4C4D2C2053";
  acc_vect( 352) <= x"10000004A44F4D4520";
  acc_vect( 353) <= x"000000000000000000";
  acc_vect( 354) <= x"11F0007B504F4D4520";
  acc_vect( 355) <= x"10000004A853545249";
  acc_vect( 356) <= x"000000000000000000";
  acc_vect( 357) <= x"11F0007B5453545249";
  acc_vect( 358) <= x"000000000000000000";
  acc_vect( 359) <= x"000000000000000000";
  acc_vect( 360) <= x"10000004804E470009";
  acc_vect( 361) <= x"000000000000000000";
  acc_vect( 362) <= x"11C0007B584E474E47";
  acc_vect( 363) <= x"000000000000000000";
  acc_vect( 364) <= x"1120007B5A00000000";
  acc_vect( 365) <= x"11F0009FB044485259";
  acc_vect( 366) <= x"11F0009FB453544F4E";
  acc_vect( 367) <= x"11F0009FB845205052";
  acc_vect( 368) <= x"11F0009FBC4F475241";
  acc_vect( 369) <= x"10000004AC4D2C2031";
  acc_vect( 370) <= x"000000000000000000";
  acc_vect( 371) <= x"11F0009FC04D2C2031";
  acc_vect( 372) <= x"10000004B027535420";
  acc_vect( 373) <= x"000000000000000000";
  acc_vect( 374) <= x"000000000000000000";
  acc_vect( 375) <= x"11F0009FC427535420";
  acc_vect( 376) <= x"11F0009FC853545249";
  acc_vect( 377) <= x"000000000000000000";
  acc_vect( 378) <= x"000000000000000000";
  acc_vect( 379) <= x"11C0009FCC4E474E47";
  acc_vect( 380) <= x"000000000000000000";
  acc_vect( 381) <= x"000000000000000000";
  acc_vect( 382) <= x"1120009FCE00000000";
  acc_vect( 383) <= x"000000000000000000";
  acc_vect( 384) <= x"10000004B40000A370";
  acc_vect( 385) <= x"000000000000000000";
  acc_vect( 386) <= x"11F000A3900000000A";
  acc_vect( 387) <= x"100000031800000384";
  acc_vect( 388) <= x"000000000000000000";
  acc_vect( 389) <= x"000000000000000000";
  acc_vect( 390) <= x"000000000000000000";
  acc_vect( 391) <= x"000000000000000000";
  acc_vect( 392) <= x"100000049044485259";
  acc_vect( 393) <= x"100000049453544F4E";
  acc_vect( 394) <= x"10000004F000000268";
  acc_vect( 395) <= x"000000000000000000";
  acc_vect( 396) <= x"000000000000000000";
  acc_vect( 397) <= x"000000000000000000";
  acc_vect( 398) <= x"000000000000000000";
  acc_vect( 399) <= x"11F0009F8000009F84";
  acc_vect( 400) <= x"000000000000000000";
  acc_vect( 401) <= x"000000000000000000";
  acc_vect( 402) <= x"10000002800000C450";
  acc_vect( 403) <= x"000000000000000000";
  acc_vect( 404) <= x"118000C45041414141";
  acc_vect( 405) <= x"000000000000000000";
  acc_vect( 406) <= x"10000002840000C520";
  acc_vect( 407) <= x"000000000000000000";
  acc_vect( 408) <= x"11F000C52000000000";
  acc_vect( 409) <= x"000000000000000000";
  acc_vect( 410) <= x"000000000000000000";
  acc_vect( 411) <= x"000000000000000000";
  acc_vect( 412) <= x"000000000000000000";
  acc_vect( 413) <= x"1000009F8000009F84";
  acc_vect( 414) <= x"10000004F40000023C";
  acc_vect( 415) <= x"000000000000000000";
  acc_vect( 416) <= x"000000000000000000";
  acc_vect( 417) <= x"000000000000000000";
  acc_vect( 418) <= x"000000000000000000";
  acc_vect( 419) <= x"11F0009F8000009F84";
  acc_vect( 420) <= x"000000000000000000";
  acc_vect( 421) <= x"100000025C0000C520";
  acc_vect( 422) <= x"10000002600000C450";
  acc_vect( 423) <= x"000000000000000000";
  acc_vect( 424) <= x"100000C45041420000";
  acc_vect( 425) <= x"000000000000000000";
  acc_vect( 426) <= x"000000000000000000";
  acc_vect( 427) <= x"000000000000000000";
  acc_vect( 428) <= x"100000C52000000000";
  acc_vect( 429) <= x"000000000000000000";
  acc_vect( 430) <= x"000000000000000000";
  acc_vect( 431) <= x"11F000C52000000001";
  acc_vect( 432) <= x"000000000000000000";
  acc_vect( 433) <= x"10000002640000C451";
  acc_vect( 434) <= x"000000000000000000";
  acc_vect( 435) <= x"114000C45142424242";
  acc_vect( 436) <= x"000000000000000000";
  acc_vect( 437) <= x"000000000000000000";
  acc_vect( 438) <= x"000000000000000000";
  acc_vect( 439) <= x"000000000000000000";
  acc_vect( 440) <= x"1000009F8000009F84";
  acc_vect( 441) <= x"000000000000000000";
  acc_vect( 442) <= x"11F0009FD800000002";
  acc_vect( 443) <= x"11F0009F9044485259";
  acc_vect( 444) <= x"11F0009F9453544F4E";
  acc_vect( 445) <= x"100000049845205052";
  acc_vect( 446) <= x"000000000000000000";
  acc_vect( 447) <= x"11F0009F9845205052";
  acc_vect( 448) <= x"100000049C4F475241";
  acc_vect( 449) <= x"000000000000000000";
  acc_vect( 450) <= x"11F0009F9C4F475241";
  acc_vect( 451) <= x"10000004F84D2C2032";
  acc_vect( 452) <= x"000000000000000000";
  acc_vect( 453) <= x"11F0009FA04D2C2032";
  acc_vect( 454) <= x"10000004FC274E4420";
  acc_vect( 455) <= x"000000000000000000";
  acc_vect( 456) <= x"11F0009FA4274E4420";
  acc_vect( 457) <= x"10000004A853545249";
  acc_vect( 458) <= x"000000000000000000";
  acc_vect( 459) <= x"11F0009FA853545249";
  acc_vect( 460) <= x"10000004804E470009";
  acc_vect( 461) <= x"000000000000000000";
  acc_vect( 462) <= x"000000000000000000";
  acc_vect( 463) <= x"11C0009FAC4E474E47";
  acc_vect( 464) <= x"000000000000000000";
  acc_vect( 465) <= x"000000000000000000";
  acc_vect( 466) <= x"1120009FAE00000000";
  acc_vect( 467) <= x"000000000000000000";
  acc_vect( 468) <= x"11F0009FD000000001";
  acc_vect( 469) <= x"000000000000000000";
  acc_vect( 470) <= x"000000000000000000";
  acc_vect( 471) <= x"000000000000000000";
  acc_vect( 472) <= x"100000050000000944";
  acc_vect( 473) <= x"000000000000000000";
  acc_vect( 474) <= x"000000000000000000";
  acc_vect( 475) <= x"000000000000000000";
  acc_vect( 476) <= x"000000000000000000";
  acc_vect( 477) <= x"11F0009F8000009F9C";
  acc_vect( 478) <= x"11F0009F7C00000002";
  acc_vect( 479) <= x"11F0009F7800000000";
  acc_vect( 480) <= x"11F0009F7400000000";
  acc_vect( 481) <= x"11F0009F7044485259";
  acc_vect( 482) <= x"11F0009F6C00009F84";
  acc_vect( 483) <= x"11F0009F68000003CE";
  acc_vect( 484) <= x"000000000000000000";
  acc_vect( 485) <= x"000000000000000000";
  acc_vect( 486) <= x"000000000000000000";
  acc_vect( 487) <= x"000000000000000000";
  acc_vect( 488) <= x"10000009A400000924";
  acc_vect( 489) <= x"000000000000000000";
  acc_vect( 490) <= x"000000000000000000";
  acc_vect( 491) <= x"000000000000000000";
  acc_vect( 492) <= x"000000000000000000";
  acc_vect( 493) <= x"000000000000000000";
  acc_vect( 494) <= x"1000009FB200005259";
  acc_vect( 495) <= x"000000000000000000";
  acc_vect( 496) <= x"000000000000000000";
  acc_vect( 497) <= x"1000009F9300000059";
  acc_vect( 498) <= x"11F0009F6400009F68";
  acc_vect( 499) <= x"000000000000000000";
  acc_vect( 500) <= x"000000000000000000";
  acc_vect( 501) <= x"000000000000000000";
  acc_vect( 502) <= x"000000000000000000";
  acc_vect( 503) <= x"000000000000000000";
  acc_vect( 504) <= x"000000000000000000";
  acc_vect( 505) <= x"000000000000000000";
  acc_vect( 506) <= x"000000000000000000";
  acc_vect( 507) <= x"000000000000000000";
  acc_vect( 508) <= x"000000000000000000";
  acc_vect( 509) <= x"000000000000000000";
  acc_vect( 510) <= x"1000009F6400009F68";
  acc_vect( 511) <= x"000000000000000000";
  acc_vect( 512) <= x"000000000000000000";
  acc_vect( 513) <= x"000000000000000000";
  acc_vect( 514) <= x"000000000000000000";
  acc_vect( 515) <= x"000000000000000000";
  acc_vect( 516) <= x"000000000000000000";
  acc_vect( 517) <= x"000000000000000000";
  acc_vect( 518) <= x"10000009A800002D14";
  acc_vect( 519) <= x"000000000000000000";
  acc_vect( 520) <= x"000000000000000000";
  acc_vect( 521) <= x"000000000000000000";
  acc_vect( 522) <= x"000000000000000000";
  acc_vect( 523) <= x"11F0009F6400009F68";
  acc_vect( 524) <= x"000000000000000000";
  acc_vect( 525) <= x"000000000000000000";
  acc_vect( 526) <= x"1000009FB044485259";
  acc_vect( 527) <= x"000000000000000000";
  acc_vect( 528) <= x"1000009F9044485259";
  acc_vect( 529) <= x"000000000000000000";
  acc_vect( 530) <= x"000000000000000000";
  acc_vect( 531) <= x"000000000000000000";
  acc_vect( 532) <= x"000000000000000000";
  acc_vect( 533) <= x"000000000000000000";
  acc_vect( 534) <= x"000000000000000000";
  acc_vect( 535) <= x"000000000000000000";
  acc_vect( 536) <= x"000000000000000000";
  acc_vect( 537) <= x"000000000000000000";
  acc_vect( 538) <= x"000000000000000000";
  acc_vect( 539) <= x"1000009FB100480000";
  acc_vect( 540) <= x"000000000000000000";
  acc_vect( 541) <= x"1000009F9100480000";
  acc_vect( 542) <= x"000000000000000000";
  acc_vect( 543) <= x"000000000000000000";
  acc_vect( 544) <= x"000000000000000000";
  acc_vect( 545) <= x"000000000000000000";
  acc_vect( 546) <= x"000000000000000000";
  acc_vect( 547) <= x"000000000000000000";
  acc_vect( 548) <= x"000000000000000000";
  acc_vect( 549) <= x"000000000000000000";
  acc_vect( 550) <= x"000000000000000000";
  acc_vect( 551) <= x"000000000000000000";
  acc_vect( 552) <= x"1000009FB200005259";
  acc_vect( 553) <= x"000000000000000000";
  acc_vect( 554) <= x"1000009F9200005259";
  acc_vect( 555) <= x"000000000000000000";
  acc_vect( 556) <= x"000000000000000000";
  acc_vect( 557) <= x"000000000000000000";
  acc_vect( 558) <= x"000000000000000000";
  acc_vect( 559) <= x"000000000000000000";
  acc_vect( 560) <= x"000000000000000000";
  acc_vect( 561) <= x"000000000000000000";
  acc_vect( 562) <= x"000000000000000000";
  acc_vect( 563) <= x"000000000000000000";
  acc_vect( 564) <= x"000000000000000000";
  acc_vect( 565) <= x"1000009FB300000059";
  acc_vect( 566) <= x"000000000000000000";
  acc_vect( 567) <= x"1000009F9300000059";
  acc_vect( 568) <= x"000000000000000000";
  acc_vect( 569) <= x"000000000000000000";
  acc_vect( 570) <= x"000000000000000000";
  acc_vect( 571) <= x"000000000000000000";
  acc_vect( 572) <= x"000000000000000000";
  acc_vect( 573) <= x"000000000000000000";
  acc_vect( 574) <= x"000000000000000000";
  acc_vect( 575) <= x"000000000000000000";
  acc_vect( 576) <= x"000000000000000000";
  acc_vect( 577) <= x"000000000000000000";
  acc_vect( 578) <= x"1000009FB453544F4E";
  acc_vect( 579) <= x"000000000000000000";
  acc_vect( 580) <= x"1000009F9453544F4E";
  acc_vect( 581) <= x"000000000000000000";
  acc_vect( 582) <= x"000000000000000000";
  acc_vect( 583) <= x"000000000000000000";
  acc_vect( 584) <= x"000000000000000000";
  acc_vect( 585) <= x"000000000000000000";
  acc_vect( 586) <= x"000000000000000000";
  acc_vect( 587) <= x"000000000000000000";
  acc_vect( 588) <= x"000000000000000000";
  acc_vect( 589) <= x"000000000000000000";
  acc_vect( 590) <= x"000000000000000000";
  acc_vect( 591) <= x"1000009FB500540000";
  acc_vect( 592) <= x"000000000000000000";
  acc_vect( 593) <= x"1000009F9500540000";
  acc_vect( 594) <= x"000000000000000000";
  acc_vect( 595) <= x"000000000000000000";
  acc_vect( 596) <= x"000000000000000000";
  acc_vect( 597) <= x"000000000000000000";
  acc_vect( 598) <= x"000000000000000000";
  acc_vect( 599) <= x"000000000000000000";
  acc_vect( 600) <= x"000000000000000000";
  acc_vect( 601) <= x"000000000000000000";
  acc_vect( 602) <= x"000000000000000000";
  acc_vect( 603) <= x"000000000000000000";
  acc_vect( 604) <= x"1000009FB600004F4E";
  acc_vect( 605) <= x"000000000000000000";
  acc_vect( 606) <= x"1000009F9600004F4E";
  acc_vect( 607) <= x"000000000000000000";
  acc_vect( 608) <= x"000000000000000000";
  acc_vect( 609) <= x"000000000000000000";
  acc_vect( 610) <= x"000000000000000000";
  acc_vect( 611) <= x"000000000000000000";
  acc_vect( 612) <= x"000000000000000000";
  acc_vect( 613) <= x"000000000000000000";
  acc_vect( 614) <= x"000000000000000000";
  acc_vect( 615) <= x"000000000000000000";
  acc_vect( 616) <= x"000000000000000000";
  acc_vect( 617) <= x"1000009FB70000004E";
  acc_vect( 618) <= x"000000000000000000";
  acc_vect( 619) <= x"1000009F970000004E";
  acc_vect( 620) <= x"000000000000000000";
  acc_vect( 621) <= x"000000000000000000";
  acc_vect( 622) <= x"000000000000000000";
  acc_vect( 623) <= x"000000000000000000";
  acc_vect( 624) <= x"000000000000000000";
  acc_vect( 625) <= x"000000000000000000";
  acc_vect( 626) <= x"000000000000000000";
  acc_vect( 627) <= x"000000000000000000";
  acc_vect( 628) <= x"000000000000000000";
  acc_vect( 629) <= x"000000000000000000";
  acc_vect( 630) <= x"1000009FB845205052";
  acc_vect( 631) <= x"000000000000000000";
  acc_vect( 632) <= x"1000009F9845205052";
  acc_vect( 633) <= x"000000000000000000";
  acc_vect( 634) <= x"000000000000000000";
  acc_vect( 635) <= x"000000000000000000";
  acc_vect( 636) <= x"000000000000000000";
  acc_vect( 637) <= x"000000000000000000";
  acc_vect( 638) <= x"000000000000000000";
  acc_vect( 639) <= x"000000000000000000";
  acc_vect( 640) <= x"000000000000000000";
  acc_vect( 641) <= x"000000000000000000";
  acc_vect( 642) <= x"000000000000000000";
  acc_vect( 643) <= x"1000009FB900200000";
  acc_vect( 644) <= x"000000000000000000";
  acc_vect( 645) <= x"1000009F9900200000";
  acc_vect( 646) <= x"000000000000000000";
  acc_vect( 647) <= x"000000000000000000";
  acc_vect( 648) <= x"000000000000000000";
  acc_vect( 649) <= x"000000000000000000";
  acc_vect( 650) <= x"000000000000000000";
  acc_vect( 651) <= x"000000000000000000";
  acc_vect( 652) <= x"000000000000000000";
  acc_vect( 653) <= x"000000000000000000";
  acc_vect( 654) <= x"000000000000000000";
  acc_vect( 655) <= x"000000000000000000";
  acc_vect( 656) <= x"1000009FBA00005052";
  acc_vect( 657) <= x"000000000000000000";
  acc_vect( 658) <= x"1000009F9A00005052";
  acc_vect( 659) <= x"000000000000000000";
  acc_vect( 660) <= x"000000000000000000";
  acc_vect( 661) <= x"000000000000000000";
  acc_vect( 662) <= x"000000000000000000";
  acc_vect( 663) <= x"000000000000000000";
  acc_vect( 664) <= x"000000000000000000";
  acc_vect( 665) <= x"000000000000000000";
  acc_vect( 666) <= x"000000000000000000";
  acc_vect( 667) <= x"000000000000000000";
  acc_vect( 668) <= x"000000000000000000";
  acc_vect( 669) <= x"1000009FBB00000052";
  acc_vect( 670) <= x"000000000000000000";
  acc_vect( 671) <= x"1000009F9B00000052";
  acc_vect( 672) <= x"000000000000000000";
  acc_vect( 673) <= x"000000000000000000";
  acc_vect( 674) <= x"000000000000000000";
  acc_vect( 675) <= x"000000000000000000";
  acc_vect( 676) <= x"000000000000000000";
  acc_vect( 677) <= x"000000000000000000";
  acc_vect( 678) <= x"000000000000000000";
  acc_vect( 679) <= x"000000000000000000";
  acc_vect( 680) <= x"000000000000000000";
  acc_vect( 681) <= x"000000000000000000";
  acc_vect( 682) <= x"1000009FBC4F475241";
  acc_vect( 683) <= x"000000000000000000";
  acc_vect( 684) <= x"1000009F9C4F475241";
  acc_vect( 685) <= x"000000000000000000";
  acc_vect( 686) <= x"000000000000000000";
  acc_vect( 687) <= x"000000000000000000";
  acc_vect( 688) <= x"000000000000000000";
  acc_vect( 689) <= x"000000000000000000";
  acc_vect( 690) <= x"000000000000000000";
  acc_vect( 691) <= x"000000000000000000";
  acc_vect( 692) <= x"000000000000000000";
  acc_vect( 693) <= x"000000000000000000";
  acc_vect( 694) <= x"000000000000000000";
  acc_vect( 695) <= x"1000009FBD00470000";
  acc_vect( 696) <= x"000000000000000000";
  acc_vect( 697) <= x"1000009F9D00470000";
  acc_vect( 698) <= x"000000000000000000";
  acc_vect( 699) <= x"000000000000000000";
  acc_vect( 700) <= x"000000000000000000";
  acc_vect( 701) <= x"000000000000000000";
  acc_vect( 702) <= x"000000000000000000";
  acc_vect( 703) <= x"000000000000000000";
  acc_vect( 704) <= x"000000000000000000";
  acc_vect( 705) <= x"000000000000000000";
  acc_vect( 706) <= x"000000000000000000";
  acc_vect( 707) <= x"000000000000000000";
  acc_vect( 708) <= x"1000009FBE00005241";
  acc_vect( 709) <= x"000000000000000000";
  acc_vect( 710) <= x"1000009F9E00005241";
  acc_vect( 711) <= x"000000000000000000";
  acc_vect( 712) <= x"000000000000000000";
  acc_vect( 713) <= x"000000000000000000";
  acc_vect( 714) <= x"000000000000000000";
  acc_vect( 715) <= x"000000000000000000";
  acc_vect( 716) <= x"000000000000000000";
  acc_vect( 717) <= x"000000000000000000";
  acc_vect( 718) <= x"000000000000000000";
  acc_vect( 719) <= x"000000000000000000";
  acc_vect( 720) <= x"000000000000000000";
  acc_vect( 721) <= x"1000009FBF00000041";
  acc_vect( 722) <= x"000000000000000000";
  acc_vect( 723) <= x"1000009F9F00000041";
  acc_vect( 724) <= x"000000000000000000";
  acc_vect( 725) <= x"000000000000000000";
  acc_vect( 726) <= x"000000000000000000";
  acc_vect( 727) <= x"000000000000000000";
  acc_vect( 728) <= x"000000000000000000";
  acc_vect( 729) <= x"000000000000000000";
  acc_vect( 730) <= x"000000000000000000";
  acc_vect( 731) <= x"000000000000000000";
  acc_vect( 732) <= x"000000000000000000";
  acc_vect( 733) <= x"000000000000000000";
  acc_vect( 734) <= x"1000009FC04D2C2031";
  acc_vect( 735) <= x"000000000000000000";
  acc_vect( 736) <= x"1000009FA04D2C2032";
  acc_vect( 737) <= x"000000000000000000";
  acc_vect( 738) <= x"000000000000000000";
  acc_vect( 739) <= x"000000000000000000";
  acc_vect( 740) <= x"000000000000000000";
  acc_vect( 741) <= x"000000000000000000";
  acc_vect( 742) <= x"000000000000000000";
  acc_vect( 743) <= x"000000000000000000";
  acc_vect( 744) <= x"000000000000000000";
  acc_vect( 745) <= x"000000000000000000";
  acc_vect( 746) <= x"000000000000000000";
  acc_vect( 747) <= x"1000009FC1002C0000";
  acc_vect( 748) <= x"000000000000000000";
  acc_vect( 749) <= x"1000009FA1002C0000";
  acc_vect( 750) <= x"000000000000000000";
  acc_vect( 751) <= x"000000000000000000";
  acc_vect( 752) <= x"000000000000000000";
  acc_vect( 753) <= x"000000000000000000";
  acc_vect( 754) <= x"000000000000000000";
  acc_vect( 755) <= x"000000000000000000";
  acc_vect( 756) <= x"000000000000000000";
  acc_vect( 757) <= x"000000000000000000";
  acc_vect( 758) <= x"000000000000000000";
  acc_vect( 759) <= x"000000000000000000";
  acc_vect( 760) <= x"1000009FC200002031";
  acc_vect( 761) <= x"000000000000000000";
  acc_vect( 762) <= x"1000009FA200002032";
  acc_vect( 763) <= x"000000000000000000";
  acc_vect( 764) <= x"000000000000000000";
  acc_vect( 765) <= x"000000000000000000";
  acc_vect( 766) <= x"000000000000000000";
  acc_vect( 767) <= x"000000000000000000";
  acc_vect( 768) <= x"000000000000000000";
  acc_vect( 769) <= x"000000000000000000";
  acc_vect( 770) <= x"000000000000000000";
  acc_vect( 771) <= x"000000000000000000";
  acc_vect( 772) <= x"000000000000000000";
  acc_vect( 773) <= x"1000009FC300000031";
  acc_vect( 774) <= x"000000000000000000";
  acc_vect( 775) <= x"1000009FA300000032";
  acc_vect( 776) <= x"000000000000000000";
  acc_vect( 777) <= x"000000000000000000";
  acc_vect( 778) <= x"000000000000000000";
  acc_vect( 779) <= x"000000000000000000";
  acc_vect( 780) <= x"000000000000000000";
  acc_vect( 781) <= x"000000000000000000";
  acc_vect( 782) <= x"000000000000000000";
  acc_vect( 783) <= x"000000000000000000";
  acc_vect( 784) <= x"000000000000000000";
  acc_vect( 785) <= x"000000000000000000";
  acc_vect( 786) <= x"000000000000000000";
  acc_vect( 787) <= x"000000000000000000";
  acc_vect( 788) <= x"1000009F6400009F68";
  acc_vect( 789) <= x"000000000000000000";
  acc_vect( 790) <= x"000000000000000000";
  acc_vect( 791) <= x"000000000000000000";
  acc_vect( 792) <= x"000000000000000000";
  acc_vect( 793) <= x"000000000000000000";
  acc_vect( 794) <= x"000000000000000000";
  acc_vect( 795) <= x"1000009F68000003CE";
  acc_vect( 796) <= x"000000000000000000";
  acc_vect( 797) <= x"000000000000000000";
  acc_vect( 798) <= x"1000009F6C00009F84";
  acc_vect( 799) <= x"000000000000000000";
  acc_vect( 800) <= x"1000009F7044485259";
  acc_vect( 801) <= x"000000000000000000";
  acc_vect( 802) <= x"1000009F7400000000";
  acc_vect( 803) <= x"000000000000000000";
  acc_vect( 804) <= x"1000009F7800000000";
  acc_vect( 805) <= x"000000000000000000";
  acc_vect( 806) <= x"1000009F7C00000002";
  acc_vect( 807) <= x"000000000000000000";
  acc_vect( 808) <= x"000000000000000000";
  acc_vect( 809) <= x"000000000000000000";
  acc_vect( 810) <= x"1000009F8000009F9C";
  acc_vect( 811) <= x"000000000000000000";
  acc_vect( 812) <= x"10000005040000C520";
  acc_vect( 813) <= x"000000000000000000";
  acc_vect( 814) <= x"11F000C52000000001";
  acc_vect( 815) <= x"1000009FD800000002";
  acc_vect( 816) <= x"000000000000000000";
  acc_vect( 817) <= x"000000000000000000";
  acc_vect( 818) <= x"000000000000000000";
  acc_vect( 819) <= x"000000000000000000";
  acc_vect( 820) <= x"100000050800000894";
  acc_vect( 821) <= x"000000000000000000";
  acc_vect( 822) <= x"000000000000000000";
  acc_vect( 823) <= x"000000000000000000";
  acc_vect( 824) <= x"000000000000000000";
  acc_vect( 825) <= x"11F0009FD400000007";
  acc_vect( 826) <= x"000000000000000000";
  acc_vect( 827) <= x"000000000000000000";
  acc_vect( 828) <= x"000000000000000000";
  acc_vect( 829) <= x"000000000000000000";
  acc_vect( 830) <= x"000000000000000000";
  acc_vect( 831) <= x"000000000000000000";
  acc_vect( 832) <= x"11F0009F8000009F84";
  acc_vect( 833) <= x"000000000000000000";
  acc_vect( 834) <= x"000000000000000000";
  acc_vect( 835) <= x"000000000000000000";
  acc_vect( 836) <= x"11F0009FD400000007";
  acc_vect( 837) <= x"000000000000000000";
  acc_vect( 838) <= x"000000000000000000";
  acc_vect( 839) <= x"000000000000000000";
  acc_vect( 840) <= x"000000000000000000";
  acc_vect( 841) <= x"1000009F8000009F84";
  acc_vect( 842) <= x"1000009FD800000002";
  acc_vect( 843) <= x"000000000000000000";
  acc_vect( 844) <= x"000000000000000000";
  acc_vect( 845) <= x"000000000000000000";
  acc_vect( 846) <= x"000000000000000000";
  acc_vect( 847) <= x"11F0009FD800000003";
  acc_vect( 848) <= x"100000050C0000C458";
  acc_vect( 849) <= x"100000051000009D34";
  acc_vect( 850) <= x"000000000000000000";
  acc_vect( 851) <= x"000000000000000000";
  acc_vect( 852) <= x"1000000514000008A4";
  acc_vect( 853) <= x"000000000000000000";
  acc_vect( 854) <= x"000000000000000000";
  acc_vect( 855) <= x"000000000000000000";
  acc_vect( 856) <= x"1000009FD400000007";
  acc_vect( 857) <= x"11F0009F8000009F9C";
  acc_vect( 858) <= x"11F0009F7C00009F84";
  acc_vect( 859) <= x"000000000000000000";
  acc_vect( 860) <= x"000000000000000000";
  acc_vect( 861) <= x"000000000000000000";
  acc_vect( 862) <= x"000000000000000000";
  acc_vect( 863) <= x"000000000000000000";
  acc_vect( 864) <= x"000000000000000000";
  acc_vect( 865) <= x"000000000000000000";
  acc_vect( 866) <= x"11F000C47800000007";
  acc_vect( 867) <= x"000000000000000000";
  acc_vect( 868) <= x"000000000000000000";
  acc_vect( 869) <= x"000000000000000000";
  acc_vect( 870) <= x"000000000000000000";
  acc_vect( 871) <= x"11F000C47C00000007";
  acc_vect( 872) <= x"000000000000000000";
  acc_vect( 873) <= x"000000000000000000";
  acc_vect( 874) <= x"000000000000000000";
  acc_vect( 875) <= x"000000000000000000";
  acc_vect( 876) <= x"000000000000000000";
  acc_vect( 877) <= x"000000000000000000";
  acc_vect( 878) <= x"000000000000000000";
  acc_vect( 879) <= x"11F000C4F000000008";
  acc_vect( 880) <= x"100000091C00C80FA0";
  acc_vect( 881) <= x"000000000000000000";
  acc_vect( 882) <= x"000000000000000000";
  acc_vect( 883) <= x"000000000000000000";
  acc_vect( 884) <= x"000000000000000000";
  acc_vect( 885) <= x"000000000000000000";
  acc_vect( 886) <= x"000000000000000000";
  acc_vect( 887) <= x"000000000000000000";
  acc_vect( 888) <= x"000000000000000000";
  acc_vect( 889) <= x"000000000000000000";
  acc_vect( 890) <= x"000000000000000000";
  acc_vect( 891) <= x"000000000000000000";
  acc_vect( 892) <= x"11F000A39400000008";
  acc_vect( 893) <= x"000000000000000000";
  acc_vect( 894) <= x"000000000000000000";
  acc_vect( 895) <= x"000000000000000000";
  acc_vect( 896) <= x"000000000000000000";
  acc_vect( 897) <= x"000000000000000000";
  acc_vect( 898) <= x"11F000A39800000008";
  acc_vect( 899) <= x"000000000000000000";
  acc_vect( 900) <= x"000000000000000000";
  acc_vect( 901) <= x"000000000000000000";
  acc_vect( 902) <= x"000000000000000000";
  acc_vect( 903) <= x"100000091C00C80FA0";
  acc_vect( 904) <= x"000000000000000000";
  acc_vect( 905) <= x"000000000000000000";
  acc_vect( 906) <= x"000000000000000000";
  acc_vect( 907) <= x"000000000000000000";
  acc_vect( 908) <= x"000000000000000000";
  acc_vect( 909) <= x"000000000000000000";
  acc_vect( 910) <= x"000000000000000000";
  acc_vect( 911) <= x"000000000000000000";
  acc_vect( 912) <= x"000000000000000000";
  acc_vect( 913) <= x"000000000000000000";
  acc_vect( 914) <= x"000000000000000000";
  acc_vect( 915) <= x"100000A3900000000A";
  acc_vect( 916) <= x"000000000000000000";
  acc_vect( 917) <= x"000000000000000000";
  acc_vect( 918) <= x"11F000A3900000000A";
  acc_vect( 919) <= x"100000091E00000FA0";
  acc_vect( 920) <= x"000000000000000000";
  acc_vect( 921) <= x"000000000000000000";
  acc_vect( 922) <= x"000000000000000000";
  acc_vect( 923) <= x"100000C47800000007";
  acc_vect( 924) <= x"000000000000000000";
  acc_vect( 925) <= x"11F000B33400000007";
  acc_vect( 926) <= x"000000000000000000";
  acc_vect( 927) <= x"10000009200000C44C";
  acc_vect( 928) <= x"000000000000000000";
  acc_vect( 929) <= x"11F000C44C00000005";
  acc_vect( 930) <= x"000000000000000000";
  acc_vect( 931) <= x"000000000000000000";
  acc_vect( 932) <= x"1000009F7C00009F84";
  acc_vect( 933) <= x"000000000000000000";
  acc_vect( 934) <= x"000000000000000000";
  acc_vect( 935) <= x"000000000000000000";
  acc_vect( 936) <= x"1000009F8000009F9C";
  acc_vect( 937) <= x"100000048C0000C454";
  acc_vect( 938) <= x"100000051800000170";
  acc_vect( 939) <= x"000000000000000000";
  acc_vect( 940) <= x"000000000000000000";
  acc_vect( 941) <= x"000000000000000000";
  acc_vect( 942) <= x"100000C45400007B2C";
  acc_vect( 943) <= x"11F0009F8000009F9C";
  acc_vect( 944) <= x"11F0009F7C00000894";
  acc_vect( 945) <= x"11F0009F7800009F84";
  acc_vect( 946) <= x"11F0009F7400000414";
  acc_vect( 947) <= x"000000000000000000";
  acc_vect( 948) <= x"000000000000000000";
  acc_vect( 949) <= x"1000007B2C00007AF8";
  acc_vect( 950) <= x"100000022C0000C454";
  acc_vect( 951) <= x"000000000000000000";
  acc_vect( 952) <= x"100000C45400007B2C";
  acc_vect( 953) <= x"000000000000000000";
  acc_vect( 954) <= x"1000007B2C00007AF8";
  acc_vect( 955) <= x"000000000000000000";
  acc_vect( 956) <= x"11F0007AF800007AF8";
  acc_vect( 957) <= x"1000007B3000000000";
  acc_vect( 958) <= x"000000000000000000";
  acc_vect( 959) <= x"11F0007AFC00000000";
  acc_vect( 960) <= x"1000007B3400000002";
  acc_vect( 961) <= x"000000000000000000";
  acc_vect( 962) <= x"11F0007B0000000002";
  acc_vect( 963) <= x"1000007B3800000028";
  acc_vect( 964) <= x"000000000000000000";
  acc_vect( 965) <= x"11F0007B0400000028";
  acc_vect( 966) <= x"1000007B3C44485259";
  acc_vect( 967) <= x"000000000000000000";
  acc_vect( 968) <= x"11F0007B0844485259";
  acc_vect( 969) <= x"1000007B4053544F4E";
  acc_vect( 970) <= x"000000000000000000";
  acc_vect( 971) <= x"11F0007B0C53544F4E";
  acc_vect( 972) <= x"1000007B4445205052";
  acc_vect( 973) <= x"000000000000000000";
  acc_vect( 974) <= x"11F0007B1045205052";
  acc_vect( 975) <= x"1000007B484F475241";
  acc_vect( 976) <= x"000000000000000000";
  acc_vect( 977) <= x"11F0007B144F475241";
  acc_vect( 978) <= x"1000007B4C4D2C2053";
  acc_vect( 979) <= x"000000000000000000";
  acc_vect( 980) <= x"11F0007B184D2C2053";
  acc_vect( 981) <= x"1000007B504F4D4520";
  acc_vect( 982) <= x"000000000000000000";
  acc_vect( 983) <= x"11F0007B1C4F4D4520";
  acc_vect( 984) <= x"1000007B5453545249";
  acc_vect( 985) <= x"000000000000000000";
  acc_vect( 986) <= x"11F0007B2053545249";
  acc_vect( 987) <= x"1000007B584E470000";
  acc_vect( 988) <= x"000000000000000000";
  acc_vect( 989) <= x"11F0007B244E470000";
  acc_vect( 990) <= x"000000000000000000";
  acc_vect( 991) <= x"11F0007B3800000005";
  acc_vect( 992) <= x"11F0007B0400000005";
  acc_vect( 993) <= x"1000007B2C00007AF8";
  acc_vect( 994) <= x"000000000000000000";
  acc_vect( 995) <= x"11F0007AF800007AF8";
  acc_vect( 996) <= x"100000023000000138";
  acc_vect( 997) <= x"000000000000000000";
  acc_vect( 998) <= x"000000000000000000";
  acc_vect( 999) <= x"000000000000000000";
  acc_vect(1000) <= x"000000000000000000";
  acc_vect(1001) <= x"11F0009F7000009F74";
  acc_vect(1002) <= x"11F0009F6C000001C2";
  acc_vect(1003) <= x"10000001640000C454";
  acc_vect(1004) <= x"000000000000000000";
  acc_vect(1005) <= x"100000C45400007B2C";
  acc_vect(1006) <= x"000000000000000000";
  acc_vect(1007) <= x"000000000000000000";
  acc_vect(1008) <= x"000000000000000000";
  acc_vect(1009) <= x"000000000000000000";
  acc_vect(1010) <= x"1000007B2C00007AF8";
  acc_vect(1011) <= x"000000000000000000";
  acc_vect(1012) <= x"11F0007AF800007AF8";
  acc_vect(1013) <= x"10000001640000C454";
  acc_vect(1014) <= x"000000000000000000";
  acc_vect(1015) <= x"100000C45400007B2C";
  acc_vect(1016) <= x"000000000000000000";
  acc_vect(1017) <= x"10000001680000C44C";
  acc_vect(1018) <= x"000000000000000000";
  acc_vect(1019) <= x"100000C44C00000005";
  acc_vect(1020) <= x"100000016C00000894";
  acc_vect(1021) <= x"000000000000000000";
  acc_vect(1022) <= x"000000000000000000";
  acc_vect(1023) <= x"000000000000000000";
  acc_vect(1024) <= x"000000000000000000";
  acc_vect(1025) <= x"11F0009F6800009F6C";
  acc_vect(1026) <= x"000000000000000000";
  acc_vect(1027) <= x"000000000000000000";
  acc_vect(1028) <= x"000000000000000000";
  acc_vect(1029) <= x"11F0007B3800000028";
  acc_vect(1030) <= x"000000000000000000";
  acc_vect(1031) <= x"000000000000000000";
  acc_vect(1032) <= x"000000000000000000";
  acc_vect(1033) <= x"000000000000000000";
  acc_vect(1034) <= x"1000009F6800009F6C";
  acc_vect(1035) <= x"000000000000000000";
  acc_vect(1036) <= x"000000000000000000";
  acc_vect(1037) <= x"1000009F6C000001C2";
  acc_vect(1038) <= x"000000000000000000";
  acc_vect(1039) <= x"000000000000000000";
  acc_vect(1040) <= x"000000000000000000";
  acc_vect(1041) <= x"000000000000000000";
  acc_vect(1042) <= x"1000009F7000009F74";
  acc_vect(1043) <= x"1000007AFC00000000";
  acc_vect(1044) <= x"000000000000000000";
  acc_vect(1045) <= x"000000000000000000";
  acc_vect(1046) <= x"000000000000000000";
  acc_vect(1047) <= x"000000000000000000";
  acc_vect(1048) <= x"11F0007B0400000006";
  acc_vect(1049) <= x"1000007B3400000002";
  acc_vect(1050) <= x"000000000000000000";
  acc_vect(1051) <= x"1000000234000009C0";
  acc_vect(1052) <= x"000000000000000000";
  acc_vect(1053) <= x"000000000000000000";
  acc_vect(1054) <= x"000000000000000000";
  acc_vect(1055) <= x"000000000000000000";
  acc_vect(1056) <= x"11F0009F7000007AF8";
  acc_vect(1057) <= x"11F0009F6C00007B2C";
  acc_vect(1058) <= x"11F0009F6800009F74";
  acc_vect(1059) <= x"11F0009F64000001D6";
  acc_vect(1060) <= x"000000000000000000";
  acc_vect(1061) <= x"000000000000000000";
  acc_vect(1062) <= x"10000009F0000009B0";
  acc_vect(1063) <= x"000000000000000000";
  acc_vect(1064) <= x"000000000000000000";
  acc_vect(1065) <= x"000000000000000000";
  acc_vect(1066) <= x"000000000000000000";
  acc_vect(1067) <= x"11F0009F6000009F64";
  acc_vect(1068) <= x"000000000000000000";
  acc_vect(1069) <= x"000000000000000000";
  acc_vect(1070) <= x"000000000000000000";
  acc_vect(1071) <= x"000000000000000000";
  acc_vect(1072) <= x"000000000000000000";
  acc_vect(1073) <= x"000000000000000000";
  acc_vect(1074) <= x"000000000000000000";
  acc_vect(1075) <= x"000000000000000000";
  acc_vect(1076) <= x"1000009F6000009F64";
  acc_vect(1077) <= x"000000000000000000";
  acc_vect(1078) <= x"000000000000000000";
  acc_vect(1079) <= x"000000000000000000";
  acc_vect(1080) <= x"000000000000000000";
  acc_vect(1081) <= x"000000000000000000";
  acc_vect(1082) <= x"11F0007B0000000002";
  acc_vect(1083) <= x"000000000000000000";
  acc_vect(1084) <= x"000000000000000000";
  acc_vect(1085) <= x"000000000000000000";
  acc_vect(1086) <= x"000000000000000000";
  acc_vect(1087) <= x"000000000000000000";
  acc_vect(1088) <= x"10000009F600002630";
  acc_vect(1089) <= x"000000000000000000";
  acc_vect(1090) <= x"000000000000000000";
  acc_vect(1091) <= x"000000000000000000";
  acc_vect(1092) <= x"000000000000000000";
  acc_vect(1093) <= x"000000000000000000";
  acc_vect(1094) <= x"000000000000000000";
  acc_vect(1095) <= x"000000000000000000";
  acc_vect(1096) <= x"11F0007B0000000001";
  acc_vect(1097) <= x"000000000000000000";
  acc_vect(1098) <= x"1000009F64000001D6";
  acc_vect(1099) <= x"000000000000000000";
  acc_vect(1100) <= x"000000000000000000";
  acc_vect(1101) <= x"1000009F6800009F74";
  acc_vect(1102) <= x"000000000000000000";
  acc_vect(1103) <= x"1000009F6C00007B2C";
  acc_vect(1104) <= x"000000000000000000";
  acc_vect(1105) <= x"000000000000000000";
  acc_vect(1106) <= x"000000000000000000";
  acc_vect(1107) <= x"1000009F7000007AF8";
  acc_vect(1108) <= x"100000022C0000C454";
  acc_vect(1109) <= x"000000000000000000";
  acc_vect(1110) <= x"100000C45400007B2C";
  acc_vect(1111) <= x"000000000000000000";
  acc_vect(1112) <= x"1000007B2C00007AF8";
  acc_vect(1113) <= x"000000000000000000";
  acc_vect(1114) <= x"11F0007AF800007AF8";
  acc_vect(1115) <= x"1000007B0400000006";
  acc_vect(1116) <= x"000000000000000000";
  acc_vect(1117) <= x"000000000000000000";
  acc_vect(1118) <= x"100000023800000894";
  acc_vect(1119) <= x"000000000000000000";
  acc_vect(1120) <= x"000000000000000000";
  acc_vect(1121) <= x"000000000000000000";
  acc_vect(1122) <= x"000000000000000000";
  acc_vect(1123) <= x"11F0009F7000009F74";
  acc_vect(1124) <= x"000000000000000000";
  acc_vect(1125) <= x"000000000000000000";
  acc_vect(1126) <= x"000000000000000000";
  acc_vect(1127) <= x"11F0007B0400000012";
  acc_vect(1128) <= x"000000000000000000";
  acc_vect(1129) <= x"000000000000000000";
  acc_vect(1130) <= x"000000000000000000";
  acc_vect(1131) <= x"000000000000000000";
  acc_vect(1132) <= x"1000009F7000009F74";
  acc_vect(1133) <= x"000000000000000000";
  acc_vect(1134) <= x"000000000000000000";
  acc_vect(1135) <= x"000000000000000000";
  acc_vect(1136) <= x"000000000000000000";
  acc_vect(1137) <= x"1000009F7400000414";
  acc_vect(1138) <= x"000000000000000000";
  acc_vect(1139) <= x"000000000000000000";
  acc_vect(1140) <= x"1000009F7800009F84";
  acc_vect(1141) <= x"000000000000000000";
  acc_vect(1142) <= x"1000009F7C00000894";
  acc_vect(1143) <= x"000000000000000000";
  acc_vect(1144) <= x"000000000000000000";
  acc_vect(1145) <= x"000000000000000000";
  acc_vect(1146) <= x"1000009F8000009F9C";
  acc_vect(1147) <= x"100000051C0000C451";
  acc_vect(1148) <= x"000000000000000000";
  acc_vect(1149) <= x"100000C45100420000";
  acc_vect(1150) <= x"000000000000000000";
  acc_vect(1151) <= x"000000000000000000";
  acc_vect(1152) <= x"000000000000000000";
  acc_vect(1153) <= x"000000000000000000";
  acc_vect(1154) <= x"000000000000000000";
  acc_vect(1155) <= x"000000000000000000";
  acc_vect(1156) <= x"10000005204D2C2033";
  acc_vect(1157) <= x"000000000000000000";
  acc_vect(1158) <= x"100000052400000924";
  acc_vect(1159) <= x"000000000000000000";
  acc_vect(1160) <= x"000000000000000000";
  acc_vect(1161) <= x"000000000000000000";
  acc_vect(1162) <= x"000000000000000000";
  acc_vect(1163) <= x"11F0009F8000009F84";
  acc_vect(1164) <= x"000000000000000000";
  acc_vect(1165) <= x"000000000000000000";
  acc_vect(1166) <= x"000000000000000000";
  acc_vect(1167) <= x"000000000000000000";
  acc_vect(1168) <= x"000000000000000000";
  acc_vect(1169) <= x"000000000000000000";
  acc_vect(1170) <= x"000000000000000000";
  acc_vect(1171) <= x"000000000000000000";
  acc_vect(1172) <= x"000000000000000000";
  acc_vect(1173) <= x"000000000000000000";
  acc_vect(1174) <= x"000000000000000000";
  acc_vect(1175) <= x"1000009F8000009F84";
  acc_vect(1176) <= x"000000000000000000";
  acc_vect(1177) <= x"000000000000000000";
  acc_vect(1178) <= x"000000000000000000";
  acc_vect(1179) <= x"1000009FD000000001";
  acc_vect(1180) <= x"000000000000000000";
  acc_vect(1181) <= x"000000000000000000";
  acc_vect(1182) <= x"000000000000000000";
  acc_vect(1183) <= x"000000000000000000";
  acc_vect(1184) <= x"000000000000000000";
  acc_vect(1185) <= x"000000000000000000";
  acc_vect(1186) <= x"000000000000000000";
  acc_vect(1187) <= x"100000051C0000C451";
  acc_vect(1188) <= x"000000000000000000";
  acc_vect(1189) <= x"100000C45100420000";
  acc_vect(1190) <= x"000000000000000000";
  acc_vect(1191) <= x"000000000000000000";
  acc_vect(1192) <= x"000000000000000000";
  acc_vect(1193) <= x"000000000000000000";
  acc_vect(1194) <= x"000000000000000000";
  acc_vect(1195) <= x"000000000000000000";
  acc_vect(1196) <= x"100000052400000924";
  acc_vect(1197) <= x"000000000000000000";
  acc_vect(1198) <= x"000000000000000000";
  acc_vect(1199) <= x"000000000000000000";
  acc_vect(1200) <= x"000000000000000000";
  acc_vect(1201) <= x"11F0009F8000009F84";
  acc_vect(1202) <= x"000000000000000000";
  acc_vect(1203) <= x"000000000000000000";
  acc_vect(1204) <= x"000000000000000000";
  acc_vect(1205) <= x"000000000000000000";
  acc_vect(1206) <= x"000000000000000000";
  acc_vect(1207) <= x"000000000000000000";
  acc_vect(1208) <= x"000000000000000000";
  acc_vect(1209) <= x"000000000000000000";
  acc_vect(1210) <= x"000000000000000000";
  acc_vect(1211) <= x"000000000000000000";
  acc_vect(1212) <= x"000000000000000000";
  acc_vect(1213) <= x"1000009F8000009F84";
  acc_vect(1214) <= x"000000000000000000";
  acc_vect(1215) <= x"000000000000000000";
  acc_vect(1216) <= x"000000000000000000";
  acc_vect(1217) <= x"1000009FD000000001";
  acc_vect(1218) <= x"000000000000000000";
  acc_vect(1219) <= x"000000000000000000";
  acc_vect(1220) <= x"000000000000000000";
  acc_vect(1221) <= x"000000000000000000";
  acc_vect(1222) <= x"000000000000000000";
  acc_vect(1223) <= x"000000000000000000";
  acc_vect(1224) <= x"000000000000000000";
  acc_vect(1225) <= x"100000051C0000C451";
  acc_vect(1226) <= x"000000000000000000";
  acc_vect(1227) <= x"100000C45100420000";
  acc_vect(1228) <= x"000000000000000000";
  acc_vect(1229) <= x"000000000000000000";
  acc_vect(1230) <= x"000000000000000000";
  acc_vect(1231) <= x"000000000000000000";
  acc_vect(1232) <= x"000000000000000000";
  acc_vect(1233) <= x"000000000000000000";
  acc_vect(1234) <= x"000000000000000000";
  acc_vect(1235) <= x"1000009FD800000003";
  acc_vect(1236) <= x"000000000000000000";
  acc_vect(1237) <= x"000000000000000000";
  acc_vect(1238) <= x"000000000000000000";
  acc_vect(1239) <= x"000000000000000000";
  acc_vect(1240) <= x"000000000000000000";
  acc_vect(1241) <= x"000000000000000000";
  acc_vect(1242) <= x"1000009FD400000007";
  acc_vect(1243) <= x"000000000000000000";
  acc_vect(1244) <= x"100000079800001ACC";
  acc_vect(1245) <= x"000000000000000000";
  acc_vect(1246) <= x"000000000000000000";
  acc_vect(1247) <= x"000000000000000000";
  acc_vect(1248) <= x"000000000000000000";
  acc_vect(1249) <= x"11F0009F8000000009";
  acc_vect(1250) <= x"000000000000000000";
  acc_vect(1251) <= x"11F0009F7C00000007";
  acc_vect(1252) <= x"000000000000000000";
  acc_vect(1253) <= x"000000000000000000";
  acc_vect(1254) <= x"000000000000000000";
  acc_vect(1255) <= x"000000000000000000";
  acc_vect(1256) <= x"000000000000000000";
  acc_vect(1257) <= x"000000000000000000";
  acc_vect(1258) <= x"000000000000000000";
  acc_vect(1259) <= x"000000000000000000";
  acc_vect(1260) <= x"000000000000000000";
  acc_vect(1261) <= x"000000000000000000";
  acc_vect(1262) <= x"000000000000000000";
  acc_vect(1263) <= x"000000000000000000";
  acc_vect(1264) <= x"000000000000000000";
  acc_vect(1265) <= x"000000000000000000";
  acc_vect(1266) <= x"000000000000000000";
  acc_vect(1267) <= x"000000000000000000";
  acc_vect(1268) <= x"000000000000000000";
  acc_vect(1269) <= x"000000000000000000";
  acc_vect(1270) <= x"000000000000000000";
  acc_vect(1271) <= x"000000000000000000";
  acc_vect(1272) <= x"000000000000000000";
  acc_vect(1273) <= x"000000000000000000";
  acc_vect(1274) <= x"000000000000000000";
  acc_vect(1275) <= x"000000000000000000";
  acc_vect(1276) <= x"000000000000000000";
  acc_vect(1277) <= x"000000000000000000";
  acc_vect(1278) <= x"000000000000000000";
  acc_vect(1279) <= x"000000000000000000";
  acc_vect(1280) <= x"000000000000000000";
  acc_vect(1281) <= x"000000000000000000";
  acc_vect(1282) <= x"000000000000000000";
  acc_vect(1283) <= x"000000000000000000";
  acc_vect(1284) <= x"000000000000000000";
  acc_vect(1285) <= x"000000000000000000";
  acc_vect(1286) <= x"000000000000000000";
  acc_vect(1287) <= x"000000000000000000";
  acc_vect(1288) <= x"000000000000000000";
  acc_vect(1289) <= x"000000000000000000";
  acc_vect(1290) <= x"000000000000000000";
  acc_vect(1291) <= x"000000000000000000";
  acc_vect(1292) <= x"000000000000000000";
  acc_vect(1293) <= x"000000000000000000";
  acc_vect(1294) <= x"000000000000000000";
  acc_vect(1295) <= x"000000000000000000";
  acc_vect(1296) <= x"000000000000000000";
  acc_vect(1297) <= x"000000000000000000";
  acc_vect(1298) <= x"000000000000000000";
  acc_vect(1299) <= x"000000000000000000";
  acc_vect(1300) <= x"000000000000000000";
  acc_vect(1301) <= x"000000000000000000";
  acc_vect(1302) <= x"000000000000000000";
  acc_vect(1303) <= x"000000000000000000";
  acc_vect(1304) <= x"000000000000000000";
  acc_vect(1305) <= x"000000000000000000";
  acc_vect(1306) <= x"000000000000000000";
  acc_vect(1307) <= x"000000000000000000";
  acc_vect(1308) <= x"000000000000000000";
  acc_vect(1309) <= x"000000000000000000";
  acc_vect(1310) <= x"000000000000000000";
  acc_vect(1311) <= x"000000000000000000";
  acc_vect(1312) <= x"000000000000000000";
  acc_vect(1313) <= x"000000000000000000";
  acc_vect(1314) <= x"000000000000000000";
  acc_vect(1315) <= x"000000000000000000";
  acc_vect(1316) <= x"000000000000000000";
  acc_vect(1317) <= x"000000000000000000";
  acc_vect(1318) <= x"000000000000000000";
  acc_vect(1319) <= x"000000000000000000";
  acc_vect(1320) <= x"000000000000000000";
  acc_vect(1321) <= x"000000000000000000";
  acc_vect(1322) <= x"1000009F7C00000007";
  acc_vect(1323) <= x"000000000000000000";
  acc_vect(1324) <= x"000000000000000000";
  acc_vect(1325) <= x"1000009F8000000009";
  acc_vect(1326) <= x"000000000000000000";
  acc_vect(1327) <= x"000000000000000000";
  acc_vect(1328) <= x"000000000000000000";
  acc_vect(1329) <= x"11F0009FD800000001";
  acc_vect(1330) <= x"000000000000000000";
  acc_vect(1331) <= x"000000000000000000";
  acc_vect(1332) <= x"000000000000000000";
  acc_vect(1333) <= x"000000000000000000";
  acc_vect(1334) <= x"000000000000000000";
  acc_vect(1335) <= x"000000000000000000";
  acc_vect(1336) <= x"000000000000000000";
  acc_vect(1337) <= x"100000079C00000110";
  acc_vect(1338) <= x"000000000000000000";
  acc_vect(1339) <= x"000000000000000000";
  acc_vect(1340) <= x"000000000000000000";
  acc_vect(1341) <= x"000000000000000000";
  acc_vect(1342) <= x"11F0009F8000009F84";
  acc_vect(1343) <= x"000000000000000000";
  acc_vect(1344) <= x"10000001300000C450";
  acc_vect(1345) <= x"000000000000000000";
  acc_vect(1346) <= x"100000C45041420000";
  acc_vect(1347) <= x"000000000000000000";
  acc_vect(1348) <= x"000000000000000000";
  acc_vect(1349) <= x"000000000000000000";
  acc_vect(1350) <= x"1000009FD800000001";
  acc_vect(1351) <= x"10000001340000C44C";
  acc_vect(1352) <= x"000000000000000000";
  acc_vect(1353) <= x"100000C44C00000005";
  acc_vect(1354) <= x"000000000000000000";
  acc_vect(1355) <= x"000000000000000000";
  acc_vect(1356) <= x"000000000000000000";
  acc_vect(1357) <= x"11F0009FD800000005";
  acc_vect(1358) <= x"000000000000000000";
  acc_vect(1359) <= x"000000000000000000";
  acc_vect(1360) <= x"000000000000000000";
  acc_vect(1361) <= x"000000000000000000";
  acc_vect(1362) <= x"1000009F8000009F84";
  acc_vect(1363) <= x"000000000000000000";
  acc_vect(1364) <= x"1000009F8800000000";
  acc_vect(1365) <= x"000000000000000000";
  acc_vect(1366) <= x"000000000000000000";
  acc_vect(1367) <= x"000000000000000000";
  acc_vect(1368) <= x"000000000000000000";
  acc_vect(1369) <= x"000000000000000000";
  acc_vect(1370) <= x"000000000000000000";
  acc_vect(1371) <= x"10000004F000000268";

end tb;
